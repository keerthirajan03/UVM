`timescale 1ns/1ps

import uvm_pkg::*;

module tb_top;
   initial begin
      run_test ("base_test");
   end

endmodule
